CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 777 301 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 778 257 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 778 219 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 778 175 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 259 376 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 256 310 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 254 248 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 256 183 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1089 320 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1089 272 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1086 214 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1085 151 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90015e-315 0
0
6 74136~
219 937 307 0 3 22
0 4 3 2
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3536 0 0
2
5.90015e-315 0
0
6 74136~
219 937 255 0 3 22
0 6 5 4
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4597 0 0
2
5.90015e-315 0
0
6 74136~
219 935 197 0 3 22
0 8 7 6
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3835 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 552 344 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 546 286 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 547 223 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 543 156 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90015e-315 0
0
6 74136~
219 381 338 0 3 22
0 13 12 9
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3108 0 0
2
5.90015e-315 0
0
6 74136~
219 377 275 0 3 22
0 14 13 10
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4299 0 0
2
5.90015e-315 0
0
6 74136~
219 374 208 0 3 22
0 15 14 11
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9672 0 0
2
5.90015e-315 0
0
20
3 1 2 0 0 4224 0 13 9 0 0 5
970 307
1077 307
1077 346
1089 346
1089 338
1 2 3 0 0 4224 0 1 13 0 0 4
789 301
913 301
913 316
921 316
0 1 4 0 0 8192 0 0 13 4 0 5
996 255
996 287
913 287
913 298
921 298
3 1 4 0 0 4224 0 14 10 0 0 5
970 255
1076 255
1076 298
1089 298
1089 290
1 2 5 0 0 4224 0 2 14 0 0 4
790 257
913 257
913 264
921 264
0 1 6 0 0 8192 0 0 14 7 0 5
995 197
995 235
913 235
913 246
921 246
3 1 6 0 0 4224 0 15 11 0 0 5
968 197
1073 197
1073 240
1086 240
1086 232
1 2 7 0 0 4224 0 3 15 0 0 4
790 219
911 219
911 206
919 206
0 1 8 0 0 8192 0 0 15 10 0 3
893 175
893 188
919 188
1 1 8 0 0 4224 0 4 12 0 0 3
790 175
1085 175
1085 169
3 1 9 0 0 4224 0 20 16 0 0 5
414 338
540 338
540 370
552 370
552 362
3 1 10 0 0 4224 0 21 17 0 0 5
410 275
534 275
534 312
546 312
546 304
3 1 11 0 0 4224 0 22 18 0 0 5
407 208
534 208
534 249
547 249
547 241
1 2 12 0 0 4224 0 5 20 0 0 4
271 376
357 376
357 347
365 347
0 1 13 0 0 4096 0 0 20 16 0 3
353 310
353 329
365 329
1 2 13 0 0 4224 0 6 21 0 0 4
268 310
353 310
353 284
361 284
0 1 14 0 0 4096 0 0 21 18 0 3
348 248
348 266
361 266
1 2 14 0 0 4224 0 7 22 0 0 4
266 248
350 248
350 217
358 217
0 1 15 0 0 8192 0 0 22 20 0 3
333 183
333 199
358 199
1 1 15 0 0 4224 0 8 19 0 0 3
268 183
543 183
543 174
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
846 354 1027 398
856 362 1016 394
31 4-Bit Gray to Binary
Converter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
297 401 478 445
307 409 467 441
31 4-Bit Binary to Gray
Converter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
