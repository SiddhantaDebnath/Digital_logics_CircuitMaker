CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 244 236 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 189 241 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 154 263 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 125 304 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 114 615 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 149 579 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 109 566 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 141 536 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 103 513 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 137 463 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 389 20 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 140 166 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 159 142 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 132 127 0 1 11
0 24
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 161 103 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 133 91 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 159 73 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 142 61 0 1 11
0 28
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 164 38 0 1 11
0 29
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 521 262 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 459 263 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 415 264 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 374 266 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90015e-315 0
0
7 74LS194
49 321 397 0 14 29
0 15 14 13 12 11 10 9 8 7
6 5 4 3 2
0
0 0 4832 90
7 74LS194
-24 -60 25 -52
2 U2
50 -11 64 -3
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 614 67 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 575 68 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 543 68 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 513 67 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 478 69 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90015e-315 0
0
7 74LS195
138 352 118 0 14 29
0 29 28 27 26 25 24 23 22 21
20 19 18 17 16
0
0 0 4832 0
7 74LS195
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 2 3 10 9 7 6 5 4 1
11 12 13 14 15 2 3 10 9 7
6 5 4 1 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3178 0 0
2
5.90015e-315 0
0
28
14 1 2 0 0 8320 0 24 20 0 0 4
357 359
357 298
521 298
521 280
13 1 3 0 0 8320 0 24 21 0 0 4
348 359
348 289
459 289
459 281
12 1 4 0 0 8320 0 24 22 0 0 4
339 359
339 295
415 295
415 282
11 1 5 0 0 4224 0 24 23 0 0 4
330 359
330 292
374 292
374 284
1 10 6 0 0 8320 0 1 24 0 0 3
256 236
312 236
312 359
1 9 7 0 0 8320 0 2 24 0 0 5
201 241
230 241
230 351
303 351
303 359
1 8 8 0 0 4224 0 3 24 0 0 3
166 263
294 263
294 359
1 7 9 0 0 4224 0 4 24 0 0 3
137 304
285 304
285 359
1 6 10 0 0 4224 0 5 24 0 0 3
126 615
357 615
357 429
1 5 11 0 0 4224 0 6 24 0 0 3
161 579
339 579
339 423
1 4 12 0 0 4224 0 7 24 0 0 3
121 566
330 566
330 423
1 3 13 0 0 4224 0 8 24 0 0 3
153 536
312 536
312 423
1 2 14 0 0 4224 0 9 24 0 0 3
115 513
303 513
303 423
1 1 15 0 0 4224 0 10 24 0 0 3
149 463
285 463
285 423
14 1 16 0 0 4224 0 30 25 0 0 3
384 154
614 154
614 85
13 1 17 0 0 4224 0 30 26 0 0 3
384 145
575 145
575 86
12 1 18 0 0 4224 0 30 27 0 0 3
384 136
543 136
543 86
11 1 19 0 0 4224 0 30 28 0 0 3
384 127
513 127
513 85
10 1 20 0 0 4224 0 30 29 0 0 3
390 118
478 118
478 87
1 9 21 0 0 8320 0 11 30 0 0 4
401 20
406 20
406 91
390 91
1 8 22 0 0 4224 0 12 30 0 0 4
152 166
306 166
306 154
320 154
1 7 23 0 0 4224 0 13 30 0 0 4
171 142
306 142
306 145
320 145
1 6 24 0 0 4224 0 14 30 0 0 4
144 127
301 127
301 136
320 136
1 5 25 0 0 4224 0 15 30 0 0 4
173 103
306 103
306 127
320 127
1 4 26 0 0 4224 0 16 30 0 0 4
145 91
291 91
291 118
314 118
1 3 27 0 0 4224 0 17 30 0 0 4
171 73
296 73
296 109
320 109
1 2 28 0 0 4224 0 18 30 0 0 4
154 61
301 61
301 100
314 100
1 1 29 0 0 4224 0 19 30 0 0 4
176 38
306 38
306 91
320 91
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 45
415 384 662 428
422 389 654 421
45 4-Bit Bidirectional Universal
Shift Register
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
383 167 614 211
390 173 606 205
49  4-Bit Parallel In Parallel 
Out Shift Register
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
