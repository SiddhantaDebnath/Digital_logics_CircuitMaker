CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 0 30 110 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 941 47 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 945 135 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 873 316 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 5.37752e-315
0
13 Logic Switch~
5 874 348 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 5.36716e-315
0
13 Logic Switch~
5 878 378 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 5.3568e-315
0
13 Logic Switch~
5 877 406 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 5.34643e-315
0
13 Logic Switch~
5 877 433 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90015e-315 5.32571e-315
0
13 Logic Switch~
5 878 463 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90015e-315 5.30499e-315
0
13 Logic Switch~
5 879 491 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90015e-315 5.26354e-315
0
13 Logic Switch~
5 881 529 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 284 509 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 282 471 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 281 443 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 280 413 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 280 386 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 281 358 0 1 11
0 24
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 277 328 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 276 296 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1368 88 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1282 169 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1183 15 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.90015e-315 0
0
6 74136~
219 1253 105 0 3 22
0 5 3 4
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9672 0 0
2
5.90015e-315 0
0
7 Ground~
168 987 94 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
5.90015e-315 0
0
6 74LS85
106 1096 207 0 14 29
0 15 14 13 12 11 10 9 8 7
2 6 5 27 3
0
0 0 5088 90
6 74LS85
48 2 90 10
2 U2
62 -8 76 0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
6369 0 0
2
5.90015e-315 5.38788e-315
0
14 Logic Display~
6 565 35 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 526 35 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 492 37 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90015e-315 0
0
6 74LS85
106 499 187 0 14 29
0 26 25 24 23 22 21 20 19 28
29 30 18 17 16
0
0 0 5088 90
6 74LS85
48 2 90 10
2 U1
62 -8 76 0
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7678 0 0
2
5.90015e-315 0
0
27
0 1 3 0 0 8192 0 0 20 4 0 4
1185 114
1185 195
1282 195
1282 187
3 1 4 0 0 4224 0 22 19 0 0 5
1286 105
1356 105
1356 114
1368 114
1368 106
0 1 5 0 0 4096 0 0 21 5 0 4
1184 96
1184 41
1183 41
1183 33
14 2 3 0 0 8320 0 24 22 0 0 3
1130 177
1130 114
1237 114
12 1 5 0 0 8320 0 24 22 0 0 3
1112 177
1112 96
1237 96
1 10 2 0 0 12416 0 23 24 0 0 4
987 88
987 84
1076 84
1076 177
1 11 6 0 0 4224 0 1 24 0 0 3
953 47
1085 47
1085 177
1 9 7 0 0 4224 0 2 24 0 0 3
957 135
1067 135
1067 177
1 8 8 0 0 8320 0 10 24 0 0 3
893 529
1130 529
1130 241
1 7 9 0 0 8320 0 9 24 0 0 3
891 491
1121 491
1121 241
1 6 10 0 0 4224 0 8 24 0 0 3
890 463
1112 463
1112 241
1 5 11 0 0 4224 0 7 24 0 0 3
889 433
1103 433
1103 241
1 4 12 0 0 4224 0 6 24 0 0 3
889 406
1094 406
1094 241
1 3 13 0 0 4224 0 5 24 0 0 3
890 378
1085 378
1085 241
1 2 14 0 0 4224 0 4 24 0 0 3
886 348
1076 348
1076 241
1 1 15 0 0 4224 0 3 24 0 0 3
885 316
1067 316
1067 241
14 1 16 0 0 4224 0 28 25 0 0 4
533 157
533 61
565 61
565 53
13 1 17 0 0 4224 0 28 26 0 0 4
524 157
524 61
526 61
526 53
12 1 18 0 0 4224 0 28 27 0 0 4
515 157
515 63
492 63
492 55
1 8 19 0 0 8320 0 11 28 0 0 3
296 509
533 509
533 221
1 7 20 0 0 8320 0 12 28 0 0 3
294 471
524 471
524 221
1 6 21 0 0 4224 0 13 28 0 0 3
293 443
515 443
515 221
1 5 22 0 0 4224 0 14 28 0 0 3
292 413
506 413
506 221
1 4 23 0 0 4224 0 15 28 0 0 3
292 386
497 386
497 221
1 3 24 0 0 4224 0 16 28 0 0 3
293 358
488 358
488 221
1 2 25 0 0 4224 0 17 28 0 0 3
289 328
479 328
479 221
1 1 26 0 0 4224 0 18 28 0 0 3
288 296
470 296
470 221
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1169 246 1316 268
1178 254 1306 270
16 5-Bit Comparator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
290 172 437 194
299 179 427 195
16 4-Bit Comparator
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
