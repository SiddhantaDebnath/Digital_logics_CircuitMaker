CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 327 631 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 331 595 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 335 568 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 370 501 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 372 480 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 373 454 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 178 28 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 95 273 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 99 243 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 91 207 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 96 164 0 1 11
0 24
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 92 132 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 95 103 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 92 75 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 92 43 0 1 11
0 28
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 924 419 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 878 424 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 839 424 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 797 426 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 757 426 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 709 429 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 674 427 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 636 434 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90015e-315 0
0
7 74LS138
19 551 516 0 14 29
0 16 15 14 11 12 13 10 9 8
7 6 5 4 3
0
0 0 5088 0
7 74LS138
-25 -61 24 -53
2 U2
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 766 113 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 730 112 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 693 114 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90015e-315 0
0
7 Ground~
168 615 78 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
5.90015e-315 0
0
5 74148
219 493 160 0 14 29
0 20 21 22 23 24 25 26 27 28
29 17 18 19 2
0
0 0 4832 0
5 74148
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 3 2 1 13 12 11 10
15 9 7 6 14 5 4 3 2 1
13 12 11 10 15 9 7 6 14 0
65 0 0 512 1 0 0 0
1 U
961 0 0
2
5.90015e-315 0
0
27
14 1 3 0 0 4224 0 24 16 0 0 3
589 552
924 552
924 437
13 1 4 0 0 4224 0 24 17 0 0 3
589 543
878 543
878 442
12 1 5 0 0 4224 0 24 18 0 0 3
589 534
839 534
839 442
11 1 6 0 0 4224 0 24 19 0 0 3
589 525
797 525
797 444
10 1 7 0 0 4224 0 24 20 0 0 3
589 516
757 516
757 444
9 1 8 0 0 4224 0 24 21 0 0 3
589 507
709 507
709 447
8 1 9 0 0 4224 0 24 22 0 0 3
589 498
674 498
674 445
7 1 10 0 0 4224 0 24 23 0 0 3
589 489
636 489
636 452
1 4 11 0 0 4224 0 1 24 0 0 4
339 631
495 631
495 534
519 534
1 5 12 0 0 4224 0 2 24 0 0 4
343 595
500 595
500 543
513 543
1 6 13 0 0 4224 0 3 24 0 0 4
347 568
505 568
505 552
513 552
1 3 14 0 0 4224 0 4 24 0 0 4
382 501
505 501
505 507
519 507
1 2 15 0 0 4224 0 5 24 0 0 4
384 480
500 480
500 498
519 498
1 1 16 0 0 4224 0 6 24 0 0 4
385 454
505 454
505 489
519 489
14 1 2 0 0 4224 0 29 28 0 0 5
531 124
601 124
601 64
615 64
615 72
11 1 17 0 0 4224 0 29 25 0 0 3
531 169
766 169
766 131
12 1 18 0 0 4224 0 29 26 0 0 3
531 160
730 160
730 130
13 1 19 0 0 4224 0 29 27 0 0 3
531 151
693 151
693 132
1 1 20 0 0 4224 0 7 29 0 0 4
190 28
432 28
432 124
455 124
1 2 21 0 0 4224 0 8 29 0 0 4
107 273
412 273
412 142
455 142
1 3 22 0 0 4224 0 9 29 0 0 4
111 243
417 243
417 151
455 151
1 4 23 0 0 4224 0 10 29 0 0 4
103 207
422 207
422 160
455 160
1 5 24 0 0 4224 0 11 29 0 0 4
108 164
427 164
427 169
455 169
1 6 25 0 0 4224 0 12 29 0 0 4
104 132
432 132
432 178
455 178
1 7 26 0 0 4224 0 13 29 0 0 4
107 103
437 103
437 187
455 187
1 8 27 0 0 4224 0 14 29 0 0 4
104 75
442 75
442 196
455 196
1 9 28 0 0 4224 0 15 29 0 0 4
104 43
447 43
447 205
455 205
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
538 583 719 607
548 591 708 607
20 Binary-Octal Decoder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
477 225 658 249
487 233 647 249
20 Octal-Binary Encoder
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
