CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
260 0 30 200 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 458 246 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 456 201 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 457 116 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 457 92 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 463 64 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 131 287 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 130 241 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 117 165 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 117 113 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 679 160 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 640 164 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90015e-315 0
0
5 4027~
219 561 246 0 7 32
0 19 5 4 5 20 2 3
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
9998 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 688 35 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 649 37 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90015e-315 0
0
5 4027~
219 553 118 0 7 32
0 21 10 9 8 22 6 7
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3835 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 322 209 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 275 213 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90015e-315 0
0
13 SR Flip-Flop~
219 215 297 0 4 9
0 14 13 11 12
0
0 0 4704 0
4 SRFF
-14 -53 14 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9323 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 319 81 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 271 89 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90015e-315 0
0
12 D Flip-Flop~
219 211 174 0 4 9
0 18 17 15 16
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
5.90015e-315 0
0
18
6 1 2 0 0 4224 0 12 10 0 0 3
591 228
679 228
679 178
7 1 3 0 0 4224 0 12 11 0 0 3
585 210
640 210
640 182
1 3 4 0 0 4224 0 1 12 0 0 4
470 246
529 246
529 219
537 219
0 4 5 0 0 4096 0 0 12 5 0 3
511 201
511 228
537 228
1 2 5 0 0 4224 0 2 12 0 0 4
468 201
529 201
529 210
537 210
6 1 6 0 0 4224 0 15 13 0 0 3
583 100
688 100
688 53
7 1 7 0 0 4224 0 15 14 0 0 3
577 82
649 82
649 55
1 4 8 0 0 4224 0 3 15 0 0 4
469 116
521 116
521 100
529 100
1 3 9 0 0 4224 0 4 15 0 0 4
469 92
521 92
521 91
529 91
1 2 10 0 0 4224 0 5 15 0 0 4
475 64
521 64
521 82
529 82
3 1 11 0 0 4224 0 18 16 0 0 3
245 279
322 279
322 227
4 1 12 0 0 4224 0 18 17 0 0 3
239 261
275 261
275 231
1 2 13 0 0 4224 0 6 18 0 0 4
143 287
183 287
183 279
191 279
1 1 14 0 0 4224 0 7 18 0 0 4
142 241
183 241
183 261
191 261
3 1 15 0 0 4224 0 21 19 0 0 3
241 156
319 156
319 99
4 1 16 0 0 4224 0 21 20 0 0 3
235 138
271 138
271 107
1 2 17 0 0 4224 0 8 21 0 0 4
129 165
179 165
179 156
187 156
1 1 18 0 0 4224 0 9 21 0 0 4
129 113
179 113
179 138
187 138
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
545 268 644 292
550 272 638 288
11 T Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
526 129 633 153
531 133 627 149
12 JK-Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
201 306 308 330
206 310 302 326
12 SR Flip Flop
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
188 170 287 194
193 174 281 190
11 D Flip Flop
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
