CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
130 0 30 100 10
487 215 1445 688
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
0 4 0.500000 0.500000
655 311 768 408
9961490 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 545 338 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44558.5 0
0
13 Logic Switch~
5 833 192 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44558.5 0
0
13 Logic Switch~
5 834 163 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44558.5 0
0
13 Logic Switch~
5 826 64 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44558.5 0
0
13 Logic Switch~
5 825 35 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
44558.5 0
0
13 Logic Switch~
5 508 81 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5572 0 0
2
44558.5 0
0
13 Logic Switch~
5 510 48 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
44558.5 0
0
13 Logic Switch~
5 226 77 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7361 0 0
2
44558.5 0
0
13 Logic Switch~
5 226 51 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4747 0 0
2
44558.5 0
0
13 Logic Switch~
5 178 367 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
972 0 0
2
44558.5 0
0
13 Logic Switch~
5 180 337 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3472 0 0
2
44558.5 0
0
13 Logic Switch~
5 449 222 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9998 0 0
2
44558.5 0
0
13 Logic Switch~
5 450 182 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3536 0 0
2
44558.5 0
0
14 Logic Display~
6 681 324 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
44558.5 0
0
9 Inverter~
13 631 338 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3835 0 0
2
44558.5 0
0
14 Logic Display~
6 997 155 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
44558.5 0
0
6 74266~
219 913 174 0 3 22
0 6 5 4
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5616 0 0
2
44558.5 0
0
14 Logic Display~
6 980 22 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
44558.5 0
0
6 74136~
219 907 45 0 3 22
0 9 8 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
317 0 0
2
44558.5 0
0
14 Logic Display~
6 690 41 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
44558.5 0
0
9 2-In NOR~
219 616 60 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4299 0 0
2
44558.5 0
0
14 Logic Display~
6 369 45 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
44558.5 0
0
10 2-In NAND~
219 301 62 0 3 22
0 15 14 13
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7876 0 0
2
44558.5 0
0
14 Logic Display~
6 383 323 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
44558.5 0
0
8 2-In OR~
219 297 343 0 3 22
0 18 17 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9172 0 0
2
44558.5 0
0
14 Logic Display~
6 717 183 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
44558.5 0
0
9 2-In AND~
219 618 196 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3820 0 0
2
44558.5 0
0
20
2 1 2 0 0 4224 0 15 14 0 0 5
652 338
669 338
669 350
681 350
681 342
1 1 3 0 0 4224 0 1 15 0 0 2
557 338
616 338
3 1 4 0 0 4224 0 17 16 0 0 5
952 174
985 174
985 181
997 181
997 173
1 2 5 0 0 4224 0 2 17 0 0 4
845 192
889 192
889 183
897 183
1 1 6 0 0 4224 0 3 17 0 0 4
846 163
889 163
889 165
897 165
3 1 7 0 0 4224 0 19 18 0 0 3
940 45
980 45
980 40
1 2 8 0 0 4224 0 4 19 0 0 4
838 64
883 64
883 54
891 54
1 1 9 0 0 4224 0 5 19 0 0 4
837 35
883 35
883 36
891 36
3 1 10 0 0 4224 0 21 20 0 0 5
655 60
678 60
678 67
690 67
690 59
1 2 11 0 0 4224 0 6 21 0 0 4
520 81
595 81
595 69
603 69
1 1 12 0 0 4224 0 7 21 0 0 4
522 48
595 48
595 51
603 51
3 1 13 0 0 4224 0 23 22 0 0 5
328 62
357 62
357 71
369 71
369 63
1 2 14 0 0 4224 0 8 23 0 0 4
238 77
269 77
269 71
277 71
1 1 15 0 0 4224 0 9 23 0 0 4
238 51
269 51
269 53
277 53
3 1 16 0 0 4224 0 25 24 0 0 5
330 343
371 343
371 349
383 349
383 341
1 2 17 0 0 4224 0 10 25 0 0 4
190 367
276 367
276 352
284 352
1 1 18 0 0 4224 0 11 25 0 0 4
192 337
276 337
276 334
284 334
3 1 19 0 0 4224 0 27 26 0 0 5
639 196
705 196
705 209
717 209
717 201
1 2 20 0 0 4224 0 12 27 0 0 4
461 222
586 222
586 205
594 205
1 1 21 0 0 4224 0 13 27 0 0 4
462 182
586 182
586 187
594 187
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
623 351 780 375
633 359 769 375
17 NOT/Inverter Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
904 191 1005 215
914 199 994 215
10 X-NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
894 64 987 88
904 72 976 88
9 X-OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
610 77 695 101
620 85 684 101
8 NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
283 83 376 107
293 91 365 107
9 NAND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
289 367 366 391
299 375 355 391
7 OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
589 233 674 257
599 241 663 257
8 AND Gate
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
