CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 130 642 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 131 600 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
961 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 129 561 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 129 525 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3409 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 130 485 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 212 269 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
5.90015e-315 5.32571e-315
0
13 Logic Switch~
5 212 300 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3780 0 0
2
5.90015e-315 5.30499e-315
0
13 Logic Switch~
5 215 329 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
5.90015e-315 5.26354e-315
0
13 Logic Switch~
5 213 364 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 204 160 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 206 125 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 203 96 0 1 11
0 24
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 203 65 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 578 579 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90015e-315 0
0
6 74136~
219 478 599 0 3 22
0 4 3 2
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3171 0 0
2
5.90015e-315 0
0
6 74136~
219 386 556 0 3 22
0 6 5 4
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4139 0 0
2
5.90015e-315 0
0
6 74136~
219 295 520 0 3 22
0 8 7 6
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
6435 0 0
2
5.90015e-315 0
0
6 74136~
219 210 493 0 3 22
0 10 9 8
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5283 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 690 348 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.90015e-315 0
0
9 Inverter~
13 642 371 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5305 0 0
2
5.90015e-315 0
0
6 74136~
219 342 328 0 3 22
0 18 17 16
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
34 0 0
2
5.90015e-315 5.36716e-315
0
6 74136~
219 456 355 0 3 22
0 16 15 14
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
969 0 0
2
5.90015e-315 5.3568e-315
0
6 74136~
219 555 376 0 3 22
0 14 13 12
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8402 0 0
2
5.90015e-315 5.34643e-315
0
14 Logic Display~
6 678 154 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90015e-315 0
0
6 74136~
219 546 172 0 3 22
0 21 20 19
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4292 0 0
2
5.90015e-315 0
0
6 74136~
219 447 151 0 3 22
0 23 22 21
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6118 0 0
2
5.90015e-315 0
0
6 74136~
219 333 124 0 3 22
0 25 24 23
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
34 0 0
2
5.90015e-315 0
0
24
3 1 2 0 0 4224 0 15 14 0 0 5
511 599
566 599
566 605
578 605
578 597
1 2 3 0 0 4224 0 1 15 0 0 4
142 642
454 642
454 608
462 608
3 1 4 0 0 4224 0 16 15 0 0 4
419 556
454 556
454 590
462 590
1 2 5 0 0 4224 0 2 16 0 0 4
143 600
362 600
362 565
370 565
3 1 6 0 0 4224 0 17 16 0 0 4
328 520
362 520
362 547
370 547
1 2 7 0 0 4224 0 3 17 0 0 4
141 561
271 561
271 529
279 529
3 1 8 0 0 4224 0 18 17 0 0 4
243 493
271 493
271 511
279 511
1 2 9 0 0 4224 0 4 18 0 0 4
141 525
186 525
186 502
194 502
1 1 10 0 0 4224 0 5 18 0 0 4
142 485
186 485
186 484
194 484
2 1 11 0 0 4224 0 20 19 0 0 3
663 371
690 371
690 366
3 1 12 0 0 4224 0 23 20 0 0 4
588 376
619 376
619 371
627 371
1 2 13 0 0 4224 0 9 23 0 0 4
225 364
436 364
436 385
539 385
3 1 14 0 0 4224 0 22 23 0 0 4
489 355
531 355
531 367
539 367
1 2 15 0 0 12416 0 8 22 0 0 4
227 329
322 329
322 364
440 364
3 1 16 0 0 4224 0 21 22 0 0 4
375 328
432 328
432 346
440 346
1 2 17 0 0 4224 0 7 21 0 0 4
224 300
313 300
313 337
326 337
1 1 18 0 0 4224 0 6 21 0 0 4
224 269
318 269
318 319
326 319
3 1 19 0 0 4224 0 25 24 0 0 5
579 172
666 172
666 180
678 180
678 172
1 2 20 0 0 4224 0 10 25 0 0 4
216 160
427 160
427 181
530 181
3 1 21 0 0 4224 0 26 25 0 0 4
480 151
522 151
522 163
530 163
1 2 22 0 0 12416 0 11 26 0 0 4
218 125
313 125
313 160
431 160
3 1 23 0 0 4224 0 27 26 0 0 4
366 124
423 124
423 142
431 142
1 2 24 0 0 4224 0 12 27 0 0 4
215 96
304 96
304 133
317 133
1 1 25 0 0 4224 0 13 27 0 0 4
215 65
309 65
309 115
317 115
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
381 657 514 681
391 665 503 681
14 Parity Checker
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
481 300 662 324
491 308 651 324
20 Odd Parity Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
462 51 651 75
472 59 640 75
21 Even Parity Generator
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
