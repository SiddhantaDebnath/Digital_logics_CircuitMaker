CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1040 1670 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
19 E:\Software\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
133
14 Logic Display~
6 1996 1948 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L24
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5130 0 0
2
44567.8 0
0
14 Logic Display~
6 1991 1791 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L23
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
44567.8 0
0
9 2-In NOR~
219 1914 1809 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U22B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
3124 0 0
2
44567.8 0
0
9 2-In NOR~
219 1808 1808 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U22A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
3421 0 0
2
44567.8 0
0
9 2-In NOR~
219 1917 1967 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U21D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
8157 0 0
2
44567.8 0
0
9 2-In NOR~
219 1812 1967 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U21C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
5572 0 0
2
44567.8 0
0
9 2-In NOR~
219 1688 2026 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U21B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
8901 0 0
2
44567.8 0
0
9 2-In NOR~
219 1587 1994 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U21A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
7361 0 0
2
44567.8 0
0
9 2-In NOR~
219 1686 1889 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U20D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
4747 0 0
2
44567.8 0
0
9 2-In NOR~
219 1486 1937 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U20C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
972 0 0
2
44567.8 0
0
9 2-In NOR~
219 1394 1936 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U20B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
3472 0 0
2
44567.8 0
0
9 2-In NOR~
219 1283 2000 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U20A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
9998 0 0
2
44567.8 0
0
9 2-In NOR~
219 1284 1874 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U17D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
3536 0 0
2
44567.8 0
0
9 2-In NOR~
219 1184 1951 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U17C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
4597 0 0
2
44567.8 0
0
13 Logic Switch~
5 1110 2078 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V30
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3835 0 0
2
44567.8 0
0
13 Logic Switch~
5 1102 2005 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V29
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3670 0 0
2
44567.8 0
0
13 Logic Switch~
5 1096 1909 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V28
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5616 0 0
2
44567.8 0
0
14 Logic Display~
6 872 2096 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L22
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
44567.8 0
0
14 Logic Display~
6 854 1904 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L21
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
44567.8 0
0
10 2-In NAND~
219 802 2114 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3108 0 0
2
44567.8 0
0
10 2-In NAND~
219 787 1922 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
4299 0 0
2
44567.8 0
0
10 2-In NAND~
219 664 1890 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
9672 0 0
2
44567.8 0
0
10 2-In NAND~
219 676 2014 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
7876 0 0
2
44567.8 0
0
10 2-In NAND~
219 551 1992 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
6369 0 0
2
44567.8 0
0
10 2-In NAND~
219 428 1984 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
9172 0 0
2
44567.8 0
0
10 2-In NAND~
219 318 2047 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
7100 0 0
2
44567.8 0
0
10 2-In NAND~
219 316 1907 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
3820 0 0
2
44567.8 0
0
10 2-In NAND~
219 208 1999 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
7678 0 0
2
44567.8 0
0
13 Logic Switch~
5 136 2120 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
961 0 0
2
44567.8 0
0
13 Logic Switch~
5 138 2051 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3178 0 0
2
44567.8 0
0
13 Logic Switch~
5 136 1960 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3409 0 0
2
44567.8 0
0
14 Logic Display~
6 1917 168 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
44567.8 0
0
14 Logic Display~
6 2030 49 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
44567.8 0
0
9 2-In NOR~
219 1676 304 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U17B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
3780 0 0
2
44567.8 0
0
9 2-In NOR~
219 1966 67 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
9265 0 0
2
44567.8 0
0
9 2-In NOR~
219 1840 66 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U16D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
9442 0 0
2
44567.8 0
0
9 2-In NOR~
219 1848 186 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U16C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
9424 0 0
2
44567.8 0
0
9 2-In NOR~
219 1746 155 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U16B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
9968 0 0
2
44567.8 0
0
9 2-In NOR~
219 1631 121 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U16A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
9281 0 0
2
44567.8 0
0
9 2-In NOR~
219 1641 195 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
8464 0 0
2
44567.8 0
0
9 2-In NOR~
219 1517 185 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
7168 0 0
2
44567.8 0
0
9 2-In NOR~
219 1421 144 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U15B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
3171 0 0
2
44567.8 0
0
9 2-In NOR~
219 1334 281 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U15A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
4139 0 0
2
44567.8 0
0
9 2-In NOR~
219 1330 190 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U10D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
6435 0 0
2
44567.8 0
0
9 2-In NOR~
219 1327 94 0 1 22
0 0
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
5283 0 0
2
44567.8 0
0
13 Logic Switch~
5 1258 362 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6874 0 0
2
44567.8 0
0
13 Logic Switch~
5 1256 241 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5305 0 0
2
44567.8 0
0
13 Logic Switch~
5 1253 165 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
34 0 0
2
44567.8 0
0
14 Logic Display~
6 1559 1316 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
44567.8 0
0
14 Logic Display~
6 1557 1206 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
44567.8 0
0
10 2-In NAND~
219 1514 1334 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
3751 0 0
2
44567.8 0
0
10 2-In NAND~
219 1509 1224 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
4292 0 0
2
44567.8 0
0
10 2-In NAND~
219 1406 1287 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6118 0 0
2
44567.8 0
0
10 2-In NAND~
219 1405 1167 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
34 0 0
2
44567.8 0
0
10 2-In NAND~
219 1293 1232 0 1 22
0 0
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
6357 0 0
2
44567.8 0
0
13 Logic Switch~
5 1226 1296 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
319 0 0
2
44567.8 0
0
13 Logic Switch~
5 1225 1181 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3976 0 0
2
44567.8 0
0
14 Logic Display~
6 571 1608 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7634 0 0
2
44567.8 0
0
14 Logic Display~
6 546 1519 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
44567.8 0
0
8 2-In OR~
219 490 1644 0 1 22
0 0
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6748 0 0
2
44567.8 0
0
9 2-In AND~
219 409 1687 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
6901 0 0
2
44567.8 0
0
9 2-In AND~
219 423 1616 0 1 22
0 0
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
842 0 0
2
44567.8 0
0
9 Inverter~
13 336 1564 0 1 22
0 0
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U7C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
3277 0 0
2
44567.8 0
0
9 Inverter~
13 204 1680 0 1 22
0 0
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
4212 0 0
2
44567.8 0
0
6 74136~
219 440 1537 0 1 22
0 0
0
0 0 608 0
7 74LS136
-24 -24 25 -16
4 U12B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
4720 0 0
2
44567.8 0
0
6 74136~
219 206 1529 0 1 22
0 0
0
0 0 608 0
7 74LS136
-24 -24 25 -16
4 U12A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
5551 0 0
2
44567.8 0
0
13 Logic Switch~
5 124 1635 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6986 0 0
2
44567.8 0
0
13 Logic Switch~
5 121 1567 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8745 0 0
2
44567.8 0
0
13 Logic Switch~
5 122 1496 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9592 0 0
2
44567.8 0
0
13 Logic Switch~
5 751 1256 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 751 1173 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 118 1165 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
631 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 116 1089 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 113 1008 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3266 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1318 845 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1312 773 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3723 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 713 874 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 712 796 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6263 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 707 575 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 706 494 0 1 11
0 32
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 107 643 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3221 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 106 546 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3215 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 115 289 0 1 11
0 45
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7903 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 111 191 0 1 11
0 50
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7121 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 114 132 0 1 11
0 51
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 919 1275 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 918 1189 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
5.90015e-315 0
0
9 2-In AND~
219 859 1293 0 3 22
0 5 4 2
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5523 0 0
2
5.90015e-315 0
0
6 74136~
219 850 1207 0 3 22
0 5 4 3
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3330 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 483 1167 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 404 1029 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.90015e-315 0
0
8 2-In OR~
219 426 1185 0 3 22
0 8 9 7
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3685 0 0
2
5.90015e-315 0
0
9 2-In AND~
219 214 1194 0 3 22
0 11 10 9
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
7849 0 0
2
5.90015e-315 0
0
9 2-In AND~
219 354 1139 0 3 22
0 12 13 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6343 0 0
2
5.90015e-315 0
0
6 74136~
219 341 1047 0 3 22
0 13 12 6
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7376 0 0
2
5.90015e-315 0
0
6 74136~
219 199 1038 0 3 22
0 11 10 13
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9156 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1756 778 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1552 716 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 1684 796 0 3 22
0 15 15 14
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
4459 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 1577 797 0 3 22
0 17 16 15
0
0 0 608 0
6 74LS02
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3760 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 1471 837 0 3 22
0 20 19 16
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
754 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 1467 734 0 3 22
0 18 20 17
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9767 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 1385 799 0 3 22
0 18 19 20
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7978 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1024 848 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1020 781 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 970 867 0 3 22
0 23 23 21
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
659 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 966 803 0 3 22
0 24 23 22
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3800 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 870 870 0 3 22
0 27 26 23
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6792 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 870 761 0 3 22
0 25 27 24
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3701 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 785 830 0 3 22
0 25 26 27
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6316 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 936 583 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 928 506 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7988 0 0
2
5.90015e-315 0
0
9 2-In AND~
219 872 602 0 3 22
0 31 30 28
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3217 0 0
2
5.90015e-315 0
0
9 Inverter~
13 810 593 0 2 22
0 32 31
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3965 0 0
2
5.90015e-315 0
0
6 74136~
219 811 527 0 3 22
0 32 30 29
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8239 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 553 564 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 490 474 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 475 582 0 3 22
0 34 37 33
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7107 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 358 476 0 3 22
0 36 35 34
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6433 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 206 717 0 3 22
0 38 38 35
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8559 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 227 467 0 3 22
0 39 39 36
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3674 0 0
2
5.90015e-315 0
0
9 2-In NOR~
219 210 591 0 3 22
0 39 38 37
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5697 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 776 279 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 862 114 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 813 133 0 3 22
0 46 42 40
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3795 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 707 296 0 3 22
0 44 43 41
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3637 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 703 191 0 3 22
0 44 45 42
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3226 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 698 85 0 3 22
0 47 44 46
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6966 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 552 167 0 3 22
0 47 45 44
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9796 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 402 158 0 3 22
0 49 48 47
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5952 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 302 215 0 3 22
0 43 50 48
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3649 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 298 91 0 3 22
0 51 43 49
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3716 0 0
2
5.90015e-315 0
0
10 2-In NAND~
219 194 160 0 3 22
0 51 50 43
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4797 0 0
2
5.90015e-315 0
0
179
3 1 0 0 0 0 0 3 2 0 0 2
1953 1809
1991 1809
3 1 0 0 0 0 0 5 1 0 0 3
1956 1967
1996 1967
1996 1966
2 0 0 0 0 0 0 5 0 0 4 3
1904 1976
1888 1976
1888 1967
3 1 0 0 0 0 0 6 5 0 0 4
1851 1967
1888 1967
1888 1958
1904 1958
2 0 0 0 0 0 0 3 0 0 6 3
1901 1818
1889 1818
1889 1808
3 1 0 0 0 0 0 4 3 0 0 4
1847 1808
1889 1808
1889 1800
1901 1800
0 1 0 0 0 0 0 0 4 19 0 3
1362 1874
1362 1799
1795 1799
3 2 0 0 0 0 0 7 6 0 0 4
1727 2026
1772 2026
1772 1976
1799 1976
1 0 0 0 0 0 0 6 0 0 10 3
1799 1958
1772 1958
1772 1889
3 2 0 0 0 0 0 9 4 0 0 4
1725 1889
1772 1889
1772 1817
1795 1817
2 0 0 0 0 0 0 7 0 0 14 2
1675 2035
1527 2035
1 0 0 0 0 0 0 7 0 0 13 3
1675 2017
1658 2017
1658 1994
3 2 0 0 0 0 0 8 9 0 0 4
1626 1994
1658 1994
1658 1898
1673 1898
1 2 0 0 0 0 0 15 8 0 0 4
1122 2078
1527 2078
1527 2003
1574 2003
1 0 0 0 0 0 0 9 0 0 16 3
1673 1880
1558 1880
1558 1936
3 1 0 0 0 0 0 10 8 0 0 6
1525 1937
1558 1937
1558 1936
1559 1936
1559 1985
1574 1985
2 0 0 0 0 0 0 10 0 0 18 3
1473 1946
1463 1946
1463 1936
3 1 0 0 0 0 0 11 10 0 0 4
1433 1936
1463 1936
1463 1928
1473 1928
3 1 0 0 0 0 0 13 11 0 0 4
1323 1874
1362 1874
1362 1927
1381 1927
3 2 0 0 0 0 0 12 11 0 0 4
1322 2000
1361 2000
1361 1945
1381 1945
1 0 0 0 0 0 0 13 0 0 26 3
1271 1865
1147 1865
1147 1909
2 0 0 0 0 0 0 12 0 0 25 3
1270 2009
1147 2009
1147 2005
1 0 0 0 0 0 0 12 0 0 24 3
1270 1991
1242 1991
1242 1951
3 2 0 0 0 0 0 14 13 0 0 4
1223 1951
1242 1951
1242 1883
1271 1883
1 2 0 0 0 0 0 16 14 0 0 4
1114 2005
1147 2005
1147 1960
1171 1960
1 1 0 0 0 0 0 17 14 0 0 4
1108 1909
1147 1909
1147 1942
1171 1942
3 1 0 0 0 0 0 20 18 0 0 2
829 2114
872 2114
0 2 0 0 0 0 0 0 20 39 0 4
383 2047
699 2047
699 2123
778 2123
1 0 0 0 0 0 0 22 0 0 38 3
640 1881
476 1881
476 1984
3 1 0 0 0 0 0 21 19 0 0 2
814 1922
854 1922
3 1 0 0 0 0 0 22 21 0 0 4
691 1890
740 1890
740 1913
763 1913
0 1 0 0 0 0 0 0 20 33 0 3
741 2004
741 2105
778 2105
3 2 0 0 0 0 0 23 21 0 0 4
703 2014
741 2014
741 1931
763 1931
2 0 0 0 0 0 0 23 0 0 37 2
652 2023
504 2023
1 0 0 0 0 0 0 23 0 0 36 3
652 2005
613 2005
613 1943
3 2 0 0 0 0 0 24 22 0 0 4
578 1992
613 1992
613 1899
640 1899
1 2 0 0 0 0 0 29 24 0 0 4
148 2120
504 2120
504 2001
527 2001
3 1 0 0 0 0 0 25 24 0 0 4
455 1984
476 1984
476 1983
527 1983
3 2 0 0 0 0 0 26 25 0 0 4
345 2047
386 2047
386 1993
404 1993
3 1 0 0 0 0 0 27 25 0 0 4
343 1907
386 1907
386 1975
404 1975
0 1 0 0 0 0 0 0 27 46 0 3
165 1960
165 1898
292 1898
2 0 0 0 0 0 0 26 0 0 45 3
294 2056
164 2056
164 2051
1 0 0 0 0 0 0 26 0 0 44 3
294 2038
267 2038
267 1999
3 2 0 0 0 0 0 28 27 0 0 4
235 1999
267 1999
267 1916
292 1916
1 2 0 0 0 0 0 30 28 0 0 4
150 2051
164 2051
164 2008
184 2008
1 1 0 0 0 0 0 31 28 0 0 4
148 1960
165 1960
165 1990
184 1990
0 2 0 0 0 0 0 0 36 50 0 3
1802 156
1802 75
1827 75
3 1 0 0 0 0 0 35 33 0 0 2
2005 67
2030 67
3 1 0 0 0 0 0 37 32 0 0 2
1887 186
1917 186
3 1 0 0 0 0 0 38 37 0 0 6
1785 155
1802 155
1802 156
1813 156
1813 177
1835 177
3 2 0 0 0 0 0 34 38 0 0 4
1715 304
1725 304
1725 164
1733 164
3 2 0 0 0 0 0 40 37 0 0 2
1680 195
1835 195
3 1 0 0 0 0 0 39 38 0 0 4
1670 121
1705 121
1705 146
1733 146
0 2 0 0 0 0 0 0 34 55 0 3
1659 303
1659 313
1663 313
0 1 0 0 0 0 0 0 34 56 0 4
1609 303
1659 303
1659 295
1663 295
1 2 0 0 0 0 0 46 40 0 0 4
1270 362
1609 362
1609 204
1628 204
2 0 0 0 0 0 0 35 0 0 58 3
1953 76
1933 76
1933 66
3 1 0 0 0 0 0 36 35 0 0 4
1879 66
1933 66
1933 58
1953 58
0 1 0 0 0 0 0 0 36 60 0 3
1494 144
1494 57
1827 57
3 1 0 0 0 0 0 42 41 0 0 4
1460 144
1494 144
1494 176
1504 176
2 0 0 0 0 0 0 39 0 0 62 3
1618 130
1613 130
1613 121
0 1 0 0 0 0 0 0 39 63 0 5
1589 185
1589 121
1613 121
1613 112
1618 112
3 1 0 0 0 0 0 41 40 0 0 4
1556 185
1589 185
1589 186
1628 186
3 2 0 0 0 0 0 44 41 0 0 3
1369 190
1369 194
1504 194
3 2 0 0 0 0 0 43 42 0 0 4
1373 281
1389 281
1389 153
1408 153
3 1 0 0 0 0 0 45 42 0 0 4
1366 94
1388 94
1388 135
1408 135
0 1 0 0 0 0 0 0 45 68 0 3
1306 103
1306 85
1314 85
0 2 0 0 0 0 0 0 45 72 0 3
1293 165
1293 103
1314 103
2 0 0 0 0 0 0 43 0 0 70 3
1321 290
1311 290
1311 272
0 1 0 0 0 0 0 0 43 71 0 3
1293 241
1293 272
1321 272
1 2 0 0 0 0 0 47 44 0 0 4
1268 241
1293 241
1293 199
1317 199
1 1 0 0 0 0 0 48 44 0 0 4
1265 165
1293 165
1293 181
1317 181
3 1 0 0 0 0 0 52 50 0 0 2
1536 1224
1557 1224
3 1 0 0 0 0 0 51 49 0 0 2
1541 1334
1559 1334
2 0 0 0 0 0 0 51 0 0 76 3
1490 1343
1472 1343
1472 1333
0 1 0 0 0 0 0 0 51 82 0 5
1345 1232
1345 1333
1472 1333
1472 1325
1490 1325
3 2 0 0 0 0 0 53 52 0 0 4
1433 1287
1458 1287
1458 1233
1485 1233
3 1 0 0 0 0 0 54 52 0 0 4
1432 1167
1458 1167
1458 1215
1485 1215
1 0 0 0 0 0 0 54 0 0 84 3
1381 1158
1260 1158
1260 1181
2 0 0 0 0 0 0 53 0 0 83 2
1382 1296
1259 1296
1 0 0 0 0 0 0 53 0 0 82 3
1382 1278
1367 1278
1367 1232
3 2 0 0 0 0 0 55 54 0 0 4
1320 1232
1367 1232
1367 1176
1381 1176
1 2 0 0 0 0 0 56 55 0 0 4
1238 1296
1260 1296
1260 1241
1269 1241
1 1 0 0 0 0 0 57 55 0 0 4
1237 1181
1260 1181
1260 1223
1269 1223
0 2 0 0 0 0 0 0 65 93 0 3
383 1626
383 1546
424 1546
3 1 0 0 0 0 0 65 59 0 0 2
473 1537
546 1537
0 2 0 0 0 0 0 0 61 97 0 3
155 1567
155 1696
385 1696
2 1 0 0 0 0 0 64 61 0 0 4
225 1680
359 1680
359 1678
385 1678
0 1 0 0 0 0 0 0 64 98 0 3
173 1521
173 1680
189 1680
3 1 0 0 0 0 0 60 58 0 0 3
523 1644
571 1644
571 1626
3 2 0 0 0 0 0 61 60 0 0 4
430 1687
460 1687
460 1653
477 1653
3 1 0 0 0 0 0 62 60 0 0 4
444 1616
460 1616
460 1635
477 1635
1 2 0 0 0 0 0 67 62 0 0 6
136 1635
359 1635
359 1626
383 1626
383 1625
399 1625
2 1 0 0 0 0 0 63 62 0 0 3
339 1582
339 1607
399 1607
0 1 0 0 0 0 0 0 63 96 0 3
355 1529
339 1529
339 1546
3 1 0 0 0 0 0 66 65 0 0 4
239 1529
355 1529
355 1528
424 1528
1 2 0 0 0 0 0 68 66 0 0 4
133 1567
162 1567
162 1538
190 1538
1 1 0 0 0 0 0 69 66 0 0 6
134 1496
162 1496
162 1521
173 1521
173 1520
190 1520
3 1 2 0 0 4224 0 88 86 0 0 2
880 1293
919 1293
3 1 3 0 0 4224 0 89 87 0 0 2
883 1207
918 1207
2 0 4 0 0 8320 0 88 0 0 103 3
835 1302
790 1302
790 1256
0 1 5 0 0 4224 0 0 88 104 0 3
819 1198
819 1284
835 1284
1 2 4 0 0 0 0 70 89 0 0 4
763 1256
791 1256
791 1216
834 1216
1 1 5 0 0 0 0 71 89 0 0 4
763 1173
791 1173
791 1198
834 1198
3 1 6 0 0 4224 0 95 91 0 0 2
374 1047
404 1047
3 1 7 0 0 4224 0 92 90 0 0 2
459 1185
483 1185
3 1 8 0 0 8320 0 94 92 0 0 4
375 1139
383 1139
383 1176
413 1176
3 2 9 0 0 4224 0 93 92 0 0 2
235 1194
413 1194
0 2 10 0 0 4224 0 0 93 115 0 3
150 1089
150 1203
190 1203
0 1 11 0 0 4224 0 0 93 116 0 3
159 1031
159 1185
190 1185
0 2 12 0 0 4096 0 0 95 113 0 3
278 1130
278 1056
325 1056
0 2 13 0 0 4224 0 0 94 114 0 3
245 1038
245 1148
330 1148
1 1 12 0 0 8320 0 72 94 0 0 3
130 1165
130 1130
330 1130
3 1 13 0 0 0 0 96 95 0 0 2
232 1038
325 1038
1 2 10 0 0 0 0 73 96 0 0 4
128 1089
150 1089
150 1047
183 1047
1 1 11 0 0 0 0 74 96 0 0 6
125 1008
149 1008
149 1031
159 1031
159 1029
183 1029
3 1 14 0 0 4224 0 99 97 0 0 2
1723 796
1756 796
2 0 15 0 0 4096 0 99 0 0 119 3
1671 805
1655 805
1655 797
3 1 15 0 0 4224 0 100 99 0 0 4
1616 797
1655 797
1655 787
1671 787
3 2 16 0 0 12416 0 101 100 0 0 4
1510 837
1524 837
1524 806
1564 806
0 1 17 0 0 4224 0 0 100 122 0 3
1524 734
1524 788
1564 788
3 1 17 0 0 0 0 102 98 0 0 2
1506 734
1552 734
1 0 18 0 0 4224 0 102 0 0 128 3
1454 725
1351 725
1351 773
2 0 19 0 0 4224 0 101 0 0 127 3
1458 846
1352 846
1352 845
1 0 20 0 0 8192 0 101 0 0 126 3
1458 828
1436 828
1436 795
3 2 20 0 0 16512 0 103 102 0 0 6
1424 799
1436 799
1436 795
1437 795
1437 743
1454 743
1 2 19 0 0 0 0 75 103 0 0 4
1330 845
1353 845
1353 808
1372 808
1 1 18 0 0 0 0 76 103 0 0 4
1324 773
1352 773
1352 790
1372 790
3 1 21 0 0 12416 0 106 104 0 0 4
997 867
1009 867
1009 866
1024 866
3 1 22 0 0 4224 0 107 105 0 0 3
993 803
1020 803
1020 799
0 2 23 0 0 4224 0 0 107 132 0 3
922 857
922 812
942 812
1 0 23 0 0 0 0 106 0 0 133 5
946 858
922 858
922 857
921 857
921 870
3 2 23 0 0 0 0 108 106 0 0 4
897 870
921 870
921 876
946 876
3 1 24 0 0 8320 0 109 107 0 0 4
897 761
920 761
920 794
942 794
1 0 25 0 0 4224 0 109 0 0 140 3
846 752
745 752
745 796
2 0 26 0 0 4224 0 108 0 0 139 3
846 879
744 879
744 874
1 0 27 0 0 8192 0 108 0 0 138 3
846 861
829 861
829 830
3 2 27 0 0 8320 0 110 109 0 0 4
812 830
830 830
830 770
846 770
1 2 26 0 0 0 0 77 110 0 0 4
725 874
745 874
745 839
761 839
1 1 25 0 0 0 0 78 110 0 0 4
724 796
745 796
745 821
761 821
3 1 28 0 0 8320 0 113 111 0 0 3
893 602
893 601
936 601
3 1 29 0 0 4224 0 115 112 0 0 3
844 527
928 527
928 524
0 2 30 0 0 8320 0 0 113 146 0 3
760 575
760 611
848 611
2 1 31 0 0 4224 0 114 113 0 0 2
831 593
848 593
0 1 32 0 0 4224 0 0 114 147 0 3
776 518
776 593
795 593
1 2 30 0 0 0 0 79 115 0 0 4
719 575
760 575
760 536
795 536
1 1 32 0 0 0 0 80 115 0 0 4
718 494
761 494
761 518
795 518
3 1 33 0 0 4224 0 118 116 0 0 2
514 582
553 582
0 1 34 0 0 4096 0 0 118 150 0 3
433 491
433 573
462 573
3 1 34 0 0 8320 0 119 117 0 0 4
397 476
397 491
490 491
490 492
3 2 35 0 0 8320 0 120 119 0 0 4
245 717
330 717
330 485
345 485
3 1 36 0 0 4224 0 121 119 0 0 2
266 467
345 467
3 2 37 0 0 4224 0 122 118 0 0 2
249 591
462 591
0 2 38 0 0 8192 0 0 120 155 0 3
177 717
177 726
193 726
0 1 38 0 0 4224 0 0 120 158 0 5
163 643
163 717
177 717
177 708
193 708
2 0 39 0 0 4096 0 121 0 0 157 3
214 476
196 476
196 465
0 1 39 0 0 4224 0 0 121 159 0 5
163 546
163 465
196 465
196 458
214 458
1 2 38 0 0 0 0 81 122 0 0 4
119 643
163 643
163 600
197 600
1 1 39 0 0 0 0 82 122 0 0 4
118 546
163 546
163 582
197 582
3 1 40 0 0 8320 0 125 124 0 0 3
840 133
840 132
862 132
3 1 41 0 0 8320 0 126 123 0 0 3
734 296
734 297
776 297
3 2 42 0 0 8320 0 127 125 0 0 4
730 191
763 191
763 142
789 142
0 2 43 0 0 12416 0 0 126 176 0 4
247 160
239 160
239 305
683 305
1 0 44 0 0 8320 0 126 0 0 166 4
683 287
629 287
629 167
639 167
2 0 45 0 0 4096 0 127 0 0 170 2
679 200
471 200
1 0 44 0 0 0 0 127 0 0 167 3
679 182
639 182
639 167
3 2 44 0 0 0 0 129 128 0 0 4
579 167
639 167
639 94
674 94
3 1 46 0 0 8320 0 128 125 0 0 4
725 85
762 85
762 124
789 124
0 1 47 0 0 8320 0 0 128 171 0 3
468 158
468 76
674 76
1 2 45 0 0 4224 0 83 129 0 0 4
127 289
471 289
471 176
528 176
3 1 47 0 0 0 0 130 129 0 0 2
429 158
528 158
3 2 48 0 0 8320 0 131 130 0 0 4
329 215
360 215
360 167
378 167
3 1 49 0 0 8320 0 132 130 0 0 4
325 91
360 91
360 149
378 149
0 2 50 0 0 8320 0 0 131 178 0 3
149 191
149 224
278 224
0 1 51 0 0 8320 0 0 132 179 0 3
149 132
149 82
274 82
0 1 43 0 0 0 0 0 131 177 0 3
247 160
247 206
278 206
3 2 43 0 0 0 0 133 132 0 0 4
221 160
249 160
249 100
274 100
1 2 50 0 0 0 0 84 133 0 0 4
123 191
149 191
149 169
170 169
1 1 51 0 0 0 0 85 133 0 0 4
126 132
149 132
149 151
170 151
66
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
1397 1736 1666 1760
1407 1744 1655 1760
31 FULL SUBTRACTOR USING NOR LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2000 1949 2101 1973
2010 1957 2090 1973
10 DIFFERENCE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1994 1788 2063 1812
2004 1796 2052 1812
6 BORROW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1052 2060 1097 2084
1062 2068 1086 2084
3 Bin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1063 1989 1092 2013
1073 1997 1081 2013
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1058 1893 1087 1917
1068 1901 1076 1917
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
320 1828 597 1852
330 1836 586 1852
32 FULL SUBTRACTOR USING NAND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
877 1900 978 1924
887 1908 967 1924
10 DIFFERENCE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
902 2100 971 2124
912 2108 960 2124
6 BORROW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
81 2105 126 2129
91 2113 115 2129
3 Bin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
85 2036 114 2060
95 2044 103 2060
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
95 1949 124 1973
105 1957 113 1973
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
1431 7 1660 31
1441 15 1649 31
26 FULL ADDER USING NOR LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
2030 46 2099 70
2040 54 2088 70
6  Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1926 164 1971 188
1936 172 1960 188
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1206 344 1251 368
1216 352 1240 368
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1214 223 1243 247
1224 231 1232 247
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1208 148 1237 172
1218 156 1226 172
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 35
1210 1100 1511 1124
1220 1108 1500 1124
35 HALF ADDER CIRCUIT USING NAND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1566 1308 1627 1332
1576 1316 1616 1332
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1571 1199 1616 1223
1581 1207 1605 1223
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1182 1285 1211 1309
1192 1293 1200 1309
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1180 1164 1209 1188
1190 1172 1198 1188
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
700 1099 1041 1123
710 1107 1030 1123
40 HALF ADDER CIRCUIT USING XOR & AND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
229 1431 434 1455
239 1439 423 1455
23 FULL SUBTRACTOR DIAGRAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
577 1625 646 1649
587 1633 635 1649
6 BORROW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
559 1508 660 1532
569 1516 649 1532
10 DIFFERENCE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
66 1619 111 1643
76 1627 100 1643
3 Bin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
81 1545 110 1569
91 1553 99 1569
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
78 1481 107 1505
88 1489 96 1505
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
369 21 606 45
379 29 595 45
27 FULL ADDER USING NAND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
50 115 79 139
60 123 68 139
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
53 176 82 200
63 184 71 200
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
55 277 100 301
65 285 89 301
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
843 134 888 158
853 142 877 158
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
748 301 809 325
758 309 798 325
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
64 527 93 551
74 535 82 551
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
64 624 93 648
74 632 82 648
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
187 398 416 422
197 406 405 422
26 HALF ADDER USING NOR LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
500 470 561 494
510 478 550 494
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
557 570 602 594
567 578 591 594
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
665 478 694 502
675 486 683 502
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
665 560 694 584
675 568 683 584
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
938 499 1015 523
948 507 1004 523
7 d=A(+)B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
947 580 1008 604
957 588 997 604
5 b=A'B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 50
642 428 1063 452
652 436 1052 452
50 HALF SUBTRACTOR CIRCUIT USING XOR, NOT & AND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1025 776 1126 800
1035 784 1115 800
10 DIFFERANCE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1033 843 1102 867
1043 851 1091 867
6 BORROW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
668 784 697 808
678 792 686 808
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
670 860 699 884
680 868 688 884
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
728 699 1005 723
738 707 994 723
32 HALF SUBTRACTOR USING NAND LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1267 757 1296 781
1277 765 1285 781
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1271 829 1300 853
1281 837 1289 853
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1761 780 1862 804
1771 788 1851 804
10 DIFFERENCE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1562 709 1631 733
1572 717 1620 733
6 BORROW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
1377 649 1646 673
1387 657 1635 673
31 HALF SUBTRACTOR USING NOR LOGIC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
70 993 99 1017
80 1001 88 1017
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
68 1072 97 1096
78 1080 86 1096
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
61 1152 106 1176
71 1160 95 1176
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
413 1029 458 1053
423 1037 447 1053
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
487 1172 548 1196
497 1180 537 1196
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
174 947 339 971
184 955 328 971
18 FULL ADDER DIAGRAM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
704 1157 733 1181
714 1165 722 1181
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
707 1240 736 1264
717 1248 725 1264
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
935 1184 980 1208
945 1192 969 1208
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
932 1269 993 1293
942 1277 982 1293
5 Carry
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
