CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1540 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
58
13 Logic Switch~
5 1854 406 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44558.5 0
0
13 Logic Switch~
5 1854 289 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44558.5 0
0
13 Logic Switch~
5 1931 126 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44558.5 0
0
13 Logic Switch~
5 1933 89 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44558.5 0
0
13 Logic Switch~
5 1520 285 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44558.5 0
0
13 Logic Switch~
5 1505 82 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5572 0 0
2
44558.5 0
0
13 Logic Switch~
5 1506 55 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
44558.5 0
0
13 Logic Switch~
5 1130 339 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7361 0 0
2
44558.5 0
0
13 Logic Switch~
5 1122 264 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4747 0 0
2
44558.5 0
0
13 Logic Switch~
5 949 51 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
972 0 0
2
44558.5 0
0
13 Logic Switch~
5 950 17 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3472 0 0
2
44558.5 0
0
13 Logic Switch~
5 452 285 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9998 0 0
2
44558.5 0
0
13 Logic Switch~
5 453 239 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3536 0 0
2
44558.5 0
0
13 Logic Switch~
5 482 78 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
44558.5 0
0
13 Logic Switch~
5 35 319 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3835 0 0
2
44558.5 0
0
13 Logic Switch~
5 32 233 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
44558.5 0
0
13 Logic Switch~
5 74 109 0 1 11
0 48
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
44558.5 0
0
13 Logic Switch~
5 74 81 0 1 11
0 49
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
44558.5 0
0
14 Logic Display~
6 2340 318 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
44558.5 0
0
9 2-In NOR~
219 2234 340 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3108 0 0
2
44558.5 0
0
9 2-In NOR~
219 2112 386 0 3 22
0 5 6 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
4299 0 0
2
44558.5 0
0
9 2-In NOR~
219 2112 302 0 3 22
0 7 5 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
9672 0 0
2
44558.5 0
0
9 2-In NOR~
219 1959 351 0 3 22
0 7 6 5
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
7876 0 0
2
44558.5 0
0
14 Logic Display~
6 2445 29 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
44558.5 0
0
9 2-In NOR~
219 2352 49 0 3 22
0 9 10 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9172 0 0
2
44558.5 0
0
9 2-In NOR~
219 2223 28 0 3 22
0 12 11 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
7100 0 0
2
44558.5 0
0
9 2-In NOR~
219 2063 173 0 3 22
0 13 13 11
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3820 0 0
2
44558.5 0
0
9 2-In NOR~
219 2058 20 0 3 22
0 14 14 12
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
7678 0 0
2
44558.5 0
0
9 2-In NOR~
219 2061 100 0 3 22
0 14 13 10
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
961 0 0
2
44558.5 0
0
14 Logic Display~
6 1687 267 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3178 0 0
2
44558.5 0
0
9 2-In NOR~
219 1612 284 0 3 22
0 16 16 15
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3409 0 0
2
44558.5 0
0
14 Logic Display~
6 1774 45 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
44558.5 0
0
9 2-In NOR~
219 1688 63 0 3 22
0 18 18 17
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8885 0 0
2
44558.5 0
0
9 2-In NOR~
219 1580 64 0 3 22
0 20 19 18
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3780 0 0
2
44558.5 0
0
14 Logic Display~
6 1416 277 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
44558.5 0
0
9 2-In NOR~
219 1324 295 0 3 22
0 23 22 21
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9442 0 0
2
44558.5 0
0
9 2-In NOR~
219 1208 337 0 3 22
0 24 24 22
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9424 0 0
2
44558.5 0
0
9 2-In NOR~
219 1209 267 0 3 22
0 25 25 23
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9968 0 0
2
44558.5 0
0
14 Logic Display~
6 1376 56 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
44558.5 0
0
10 2-In NAND~
219 1301 71 0 3 22
0 27 28 26
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8464 0 0
2
44558.5 0
0
10 2-In NAND~
219 1219 121 0 3 22
0 30 29 28
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7168 0 0
2
44558.5 0
0
10 2-In NAND~
219 1119 157 0 3 22
0 32 32 29
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3171 0 0
2
44558.5 0
0
10 2-In NAND~
219 1118 101 0 3 22
0 31 31 30
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4139 0 0
2
44558.5 0
0
10 2-In NAND~
219 1222 32 0 3 22
0 31 32 27
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6435 0 0
2
44558.5 0
0
14 Logic Display~
6 960 217 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5283 0 0
2
44558.5 0
0
10 2-In NAND~
219 884 236 0 3 22
0 35 34 33
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6874 0 0
2
44558.5 0
0
10 2-In NAND~
219 742 281 0 3 22
0 36 37 34
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5305 0 0
2
44558.5 0
0
10 2-In NAND~
219 741 194 0 3 22
0 38 36 35
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
34 0 0
2
44558.5 0
0
10 2-In NAND~
219 582 249 0 3 22
0 38 37 36
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
969 0 0
2
44558.5 0
0
14 Logic Display~
6 652 61 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
44558.5 0
0
10 2-In NAND~
219 581 79 0 3 22
0 40 40 39
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3751 0 0
2
44558.5 0
0
14 Logic Display~
6 345 247 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
44558.5 0
0
10 2-In NAND~
219 253 265 0 3 22
0 43 42 41
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6118 0 0
2
44558.5 0
0
10 2-In NAND~
219 117 319 0 3 22
0 44 44 42
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
34 0 0
2
44558.5 0
0
10 2-In NAND~
219 116 234 0 3 22
0 45 45 43
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6357 0 0
2
44558.5 0
0
14 Logic Display~
6 348 72 0 1 2
10 46
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
319 0 0
2
44558.5 0
0
10 2-In NAND~
219 273 88 0 3 22
0 47 47 46
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3976 0 0
2
44558.5 0
0
10 2-In NAND~
219 166 90 0 3 22
0 49 48 47
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7634 0 0
2
44558.5 0
0
70
3 1 2 0 0 4224 0 20 19 0 0 3
2273 340
2340 340
2340 336
3 2 3 0 0 4224 0 21 20 0 0 4
2151 386
2213 386
2213 349
2221 349
3 1 4 0 0 4224 0 22 20 0 0 4
2151 302
2213 302
2213 331
2221 331
0 1 5 0 0 4096 0 0 21 5 0 3
2091 351
2091 377
2099 377
3 2 5 0 0 4224 0 23 22 0 0 4
1998 351
2091 351
2091 311
2099 311
0 2 6 0 0 4096 0 0 23 8 0 3
1904 406
1904 360
1946 360
0 1 7 0 0 4096 0 0 23 9 0 3
1908 289
1908 342
1946 342
1 2 6 0 0 4224 0 1 21 0 0 4
1866 406
2091 406
2091 395
2099 395
1 1 7 0 0 4224 0 2 22 0 0 4
1866 289
2091 289
2091 293
2099 293
3 1 8 0 0 4224 0 25 24 0 0 5
2391 49
2433 49
2433 55
2445 55
2445 47
3 1 9 0 0 4224 0 26 25 0 0 4
2262 28
2331 28
2331 40
2339 40
3 2 10 0 0 4224 0 29 25 0 0 4
2100 100
2331 100
2331 58
2339 58
3 2 11 0 0 8320 0 27 26 0 0 4
2102 173
2202 173
2202 37
2210 37
3 1 12 0 0 4224 0 28 26 0 0 4
2097 20
2202 20
2202 19
2210 19
0 1 13 0 0 8192 0 0 27 16 0 3
2029 182
2029 164
2050 164
0 2 13 0 0 8192 0 0 27 19 0 3
1992 126
1992 182
2050 182
0 2 14 0 0 4096 0 0 28 18 0 3
2028 11
2028 29
2045 29
0 1 14 0 0 4096 0 0 28 20 0 3
1993 89
1993 11
2045 11
1 2 13 0 0 4224 0 3 29 0 0 4
1943 126
2040 126
2040 109
2048 109
1 1 14 0 0 4224 0 4 29 0 0 4
1945 89
2040 89
2040 91
2048 91
3 1 15 0 0 4224 0 31 30 0 0 5
1651 284
1675 284
1675 293
1687 293
1687 285
0 2 16 0 0 4096 0 0 31 23 0 3
1591 285
1591 293
1599 293
1 1 16 0 0 4224 0 5 31 0 0 4
1532 285
1591 285
1591 275
1599 275
3 1 17 0 0 4224 0 33 32 0 0 5
1727 63
1762 63
1762 71
1774 71
1774 63
0 2 18 0 0 4096 0 0 33 26 0 3
1667 64
1667 72
1675 72
3 1 18 0 0 4224 0 34 33 0 0 4
1619 64
1667 64
1667 54
1675 54
1 2 19 0 0 4224 0 6 34 0 0 4
1517 82
1559 82
1559 73
1567 73
1 1 20 0 0 4224 0 7 34 0 0 2
1518 55
1567 55
3 1 21 0 0 4224 0 36 35 0 0 5
1363 295
1404 295
1404 303
1416 303
1416 295
3 2 22 0 0 4224 0 37 36 0 0 4
1247 337
1303 337
1303 304
1311 304
3 1 23 0 0 4224 0 38 36 0 0 4
1248 267
1303 267
1303 286
1311 286
0 2 24 0 0 8192 0 0 37 33 0 3
1187 339
1187 346
1195 346
1 1 24 0 0 4224 0 8 37 0 0 4
1142 339
1187 339
1187 328
1195 328
0 2 25 0 0 4096 0 0 38 35 0 3
1188 264
1188 276
1196 276
1 1 25 0 0 4224 0 9 38 0 0 4
1134 264
1188 264
1188 258
1196 258
3 1 26 0 0 4224 0 40 39 0 0 5
1328 71
1364 71
1364 82
1376 82
1376 74
3 1 27 0 0 8320 0 44 40 0 0 4
1249 32
1269 32
1269 62
1277 62
3 2 28 0 0 8320 0 41 40 0 0 4
1246 121
1269 121
1269 80
1277 80
3 2 29 0 0 4224 0 42 41 0 0 4
1146 157
1187 157
1187 130
1195 130
3 1 30 0 0 4224 0 43 41 0 0 4
1145 101
1187 101
1187 112
1195 112
0 1 31 0 0 4096 0 0 43 42 0 3
1086 110
1086 92
1094 92
0 2 31 0 0 4096 0 0 43 46 0 3
1074 17
1074 110
1094 110
0 1 32 0 0 8192 0 0 42 44 0 3
1076 166
1076 148
1095 148
0 2 32 0 0 4096 0 0 42 45 0 3
1031 51
1031 166
1095 166
1 2 32 0 0 4224 0 10 44 0 0 4
961 51
1190 51
1190 41
1198 41
1 1 31 0 0 4224 0 11 44 0 0 4
962 17
1190 17
1190 23
1198 23
3 1 33 0 0 4224 0 46 45 0 0 5
911 236
948 236
948 243
960 243
960 235
3 2 34 0 0 4224 0 47 46 0 0 4
769 281
852 281
852 245
860 245
3 1 35 0 0 4224 0 48 46 0 0 4
768 194
852 194
852 227
860 227
0 1 36 0 0 4096 0 0 47 51 0 3
707 249
707 272
718 272
3 2 36 0 0 4224 0 49 48 0 0 4
609 249
709 249
709 203
717 203
0 2 37 0 0 8320 0 0 47 54 0 3
506 285
506 290
718 290
0 1 38 0 0 8320 0 0 48 55 0 3
508 239
508 185
717 185
1 2 37 0 0 0 0 12 49 0 0 4
464 285
550 285
550 258
558 258
1 1 38 0 0 0 0 13 49 0 0 4
465 239
550 239
550 240
558 240
3 1 39 0 0 4224 0 51 50 0 0 5
608 79
640 79
640 87
652 87
652 79
0 2 40 0 0 4096 0 0 51 58 0 3
548 78
548 88
557 88
1 1 40 0 0 4224 0 14 51 0 0 4
494 78
549 78
549 70
557 70
3 1 41 0 0 4224 0 53 52 0 0 5
280 265
333 265
333 273
345 273
345 265
3 2 42 0 0 4224 0 54 53 0 0 4
144 319
221 319
221 274
229 274
3 1 43 0 0 4224 0 55 53 0 0 4
143 234
221 234
221 256
229 256
0 2 44 0 0 4096 0 0 54 63 0 3
85 319
85 328
93 328
1 1 44 0 0 4224 0 15 54 0 0 4
47 319
85 319
85 310
93 310
0 2 45 0 0 4096 0 0 55 65 0 3
84 233
84 243
92 243
1 1 45 0 0 4224 0 16 55 0 0 4
44 233
84 233
84 225
92 225
3 1 46 0 0 4224 0 57 56 0 0 5
300 88
336 88
336 98
348 98
348 90
3 2 47 0 0 4096 0 58 57 0 0 4
193 90
236 90
236 97
249 97
3 1 47 0 0 4224 0 58 57 0 0 4
193 90
241 90
241 79
249 79
1 2 48 0 0 4224 0 17 58 0 0 4
86 109
134 109
134 99
142 99
1 1 49 0 0 4224 0 18 58 0 0 2
86 81
142 81
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
1987 462 2128 486
1997 470 2117 486
15 X-NOR using NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
2001 199 2134 223
2011 207 2123 223
14 X-OR using NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1573 309 1698 333
1583 317 1687 333
13 NOT using NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1578 89 1695 113
1588 97 1684 113
12 OR using NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1193 371 1318 395
1203 379 1307 395
13 AND using NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1102 176 1251 200
1112 184 1240 200
16 X-NOR using NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
533 311 674 335
543 319 663 335
15 X-OR using NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
557 105 690 129
567 113 679 129
14 NOT using NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
81 350 206 374
91 358 195 374
13 OR using NAND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
155 115 288 139
165 123 277 139
14 AND using NAND
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
