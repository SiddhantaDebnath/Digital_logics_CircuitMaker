CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
940 0 30 150 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
54
13 Logic Switch~
5 1075 183 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V33
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6357 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1073 157 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V32
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
319 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1032 121 0 1 11
0 12
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V31
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3976 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1037 99 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V30
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7634 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1060 57 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V29
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
523 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 1061 29 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V28
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 571 431 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V27
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6901 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 572 407 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
842 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 586 357 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3277 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 585 331 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4212 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 786 103 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4720 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 790 77 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5551 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 790 51 0 1 11
0 28
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6986 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 789 26 0 1 11
0 29
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8745 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 544 250 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9592 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 544 214 0 1 11
0 31
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 543 181 0 1 11
0 32
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 541 147 0 1 11
0 33
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
631 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 541 117 0 1 11
0 34
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 541 90 0 1 11
0 35
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3266 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 539 62 0 1 11
0 36
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 538 32 0 1 11
0 37
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3723 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 150 210 0 1 11
0 50
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
3440 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 321 207 0 1 11
0 39
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6263 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 115 393 0 1 11
0 40
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 115 359 0 1 11
0 41
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 115 325 0 1 11
0 42
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3221 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 115 301 0 1 11
0 43
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3215 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 117 278 0 1 11
0 44
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7903 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 99 176 0 1 11
0 46
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7121 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 107 113 0 1 11
0 47
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 110 92 0 1 11
0 48
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 112 62 0 1 11
0 49
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7804 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1557 18 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1517 23 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1474 23 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1431 25 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1390 22 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1343 21 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1302 17 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 1265 20 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
5.90015e-315 0
0
7 74LS155
120 1189 90 0 14 29
0 15 14 13 12 11 10 9 8 7
6 5 4 3 2
0
0 0 4832 0
7 74LS155
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 13 14 15 4 5 6
7 12 11 10 9 1 2 3 13 14
15 4 5 6 7 12 11 10 9 0
65 0 0 0 1 0 0 0
1 U
9156 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 899 295 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 865 296 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 829 298 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 793 300 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
5.90015e-315 0
0
7 74LS155
120 715 385 0 14 29
0 23 22 21 20 51 52 19 18 17
16 53 54 55 56
0
0 0 4832 0
7 74LS155
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 13 14 15 4 5 6
7 12 11 10 9 1 2 3 13 14
15 4 5 6 7 12 11 10 9 0
65 0 0 512 1 0 0 0
1 U
754 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 902 98 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 857 101 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7978 0 0
2
5.90015e-315 0
0
7 74LS151
20 690 105 0 14 29
0 37 36 35 34 33 32 31 30 26
29 28 27 25 24
0
0 0 4832 0
7 74LS151
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
3142 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 395 239 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
5.90015e-315 0
0
7 74LS153
119 244 307 0 14 29
0 57 44 43 42 41 40 58 59 60
61 39 62 38 63
0
0 0 4832 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
659 0 0
2
5.90015e-315 0
0
14 Logic Display~
6 355 67 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
5.90015e-315 0
0
7 74LS157
122 243 121 0 14 29
0 49 48 47 64 65 66 67 68 69
46 45 70 71 72
0
0 0 4832 0
6 74F157
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 512 1 0 0 0
1 U
6792 0 0
2
5.90015e-315 0
0
49
1 1 0 0 0 0 0 23 52 0 0 4
162 210
204 210
204 271
212 271
14 1 2 0 0 4224 0 42 34 0 0 3
1227 126
1557 126
1557 36
13 1 3 0 0 4224 0 42 35 0 0 3
1227 117
1517 117
1517 41
12 1 4 0 0 4224 0 42 36 0 0 3
1227 108
1474 108
1474 41
11 1 5 0 0 4224 0 42 37 0 0 3
1227 99
1431 99
1431 43
10 1 6 0 0 4224 0 42 38 0 0 3
1227 90
1390 90
1390 40
9 1 7 0 0 4224 0 42 39 0 0 3
1227 81
1343 81
1343 39
8 1 8 0 0 4224 0 42 40 0 0 3
1227 72
1302 72
1302 35
7 1 9 0 0 4224 0 42 41 0 0 3
1227 63
1265 63
1265 38
1 6 10 0 0 8320 0 1 42 0 0 4
1087 183
1138 183
1138 126
1151 126
1 5 11 0 0 4224 0 2 42 0 0 4
1085 157
1143 157
1143 117
1151 117
1 4 12 0 0 4224 0 3 42 0 0 4
1044 121
1138 121
1138 99
1157 99
1 3 13 0 0 4224 0 4 42 0 0 4
1049 99
1143 99
1143 90
1157 90
1 2 14 0 0 4224 0 5 42 0 0 4
1072 57
1138 57
1138 72
1151 72
1 1 15 0 0 4224 0 6 42 0 0 4
1073 29
1143 29
1143 63
1157 63
10 1 16 0 0 4224 0 47 43 0 0 3
753 385
899 385
899 313
9 1 17 0 0 4224 0 47 44 0 0 3
753 376
865 376
865 314
8 1 18 0 0 4224 0 47 45 0 0 3
753 367
829 367
829 316
7 1 19 0 0 4224 0 47 46 0 0 3
753 358
793 358
793 318
1 4 20 0 0 4224 0 7 47 0 0 4
583 431
664 431
664 394
683 394
1 3 21 0 0 4224 0 8 47 0 0 4
584 407
669 407
669 385
683 385
1 2 22 0 0 4224 0 9 47 0 0 4
598 357
664 357
664 367
677 367
1 1 23 0 0 4224 0 10 47 0 0 4
597 331
669 331
669 358
683 358
14 1 24 0 0 4224 0 50 48 0 0 3
728 141
902 141
902 116
13 1 25 0 0 4224 0 50 49 0 0 3
722 132
857 132
857 119
1 9 26 0 0 12416 0 11 50 0 0 6
798 103
807 103
807 93
741 93
741 78
728 78
1 12 27 0 0 12416 0 12 50 0 0 6
802 77
817 77
817 114
736 114
736 105
722 105
1 11 28 0 0 12416 0 13 50 0 0 6
802 51
812 51
812 92
736 92
736 96
722 96
1 10 29 0 0 12416 0 14 50 0 0 4
801 26
808 26
808 87
722 87
1 8 30 0 0 8320 0 15 50 0 0 4
556 250
635 250
635 141
658 141
1 7 31 0 0 4224 0 16 50 0 0 4
556 214
640 214
640 132
658 132
1 6 32 0 0 4224 0 17 50 0 0 4
555 181
650 181
650 123
658 123
1 5 33 0 0 4224 0 18 50 0 0 4
553 147
645 147
645 114
658 114
1 4 34 0 0 4224 0 19 50 0 0 4
553 117
650 117
650 105
658 105
1 3 35 0 0 4224 0 20 50 0 0 4
553 90
650 90
650 96
658 96
1 2 36 0 0 4224 0 21 50 0 0 4
551 62
645 62
645 87
658 87
1 1 37 0 0 4224 0 22 50 0 0 4
550 32
650 32
650 78
658 78
13 1 38 0 0 4224 0 52 51 0 0 3
276 289
395 289
395 257
1 11 39 0 0 8320 0 24 52 0 0 4
333 207
338 207
338 271
282 271
1 6 40 0 0 8320 0 25 52 0 0 4
127 393
194 393
194 316
212 316
1 5 41 0 0 4224 0 26 52 0 0 4
127 359
204 359
204 307
212 307
1 4 42 0 0 4224 0 27 52 0 0 4
127 325
199 325
199 298
212 298
1 3 43 0 0 4224 0 28 52 0 0 4
127 301
204 301
204 289
212 289
1 2 44 0 0 4224 0 29 52 0 0 4
129 278
204 278
204 280
212 280
11 1 45 0 0 4224 0 54 53 0 0 3
275 103
355 103
355 85
1 10 46 0 0 4224 0 30 54 0 0 4
111 176
197 176
197 166
205 166
1 3 47 0 0 4224 0 31 54 0 0 4
119 113
197 113
197 103
211 103
1 2 48 0 0 4224 0 32 54 0 0 4
122 92
197 92
197 94
211 94
1 1 49 0 0 4224 0 33 54 0 0 4
124 62
197 62
197 85
211 85
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
1181 145 1364 169
1188 151 1356 167
21 1-line to 8-line DMux
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
714 441 897 465
721 446 889 462
21 1-line to 4-line DMux
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
696 157 799 181
703 163 791 179
11 8-input Mux
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
226 447 329 471
233 453 321 469
11 4-input Mux
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
223 19 326 43
230 25 318 41
11 2-input Mux
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
