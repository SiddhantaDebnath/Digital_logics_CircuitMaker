CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 460 30 150 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
22 D:\Digital Lab\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 303 233 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 337 198 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 284 171 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 645 133 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 589 149 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 545 179 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90015e-315 0
0
13 Logic Switch~
5 399 707 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44567.5 0
0
13 Logic Switch~
5 399 682 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44567.5 1
0
13 Logic Switch~
5 400 657 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44567.5 2
0
13 Logic Switch~
5 353 443 0 1 11
0 26
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44567.5 3
0
13 Logic Switch~
5 354 416 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44567.5 4
0
13 Logic Switch~
5 372 392 0 1 11
0 28
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44567.5 5
0
13 Logic Switch~
5 347 347 0 1 11
0 29
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
44567.5 6
0
13 Logic Switch~
5 353 320 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
44567.5 7
0
13 Logic Switch~
5 412 304 0 1 11
0 31
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
44567.5 8
0
13 Logic Switch~
5 414 285 0 1 11
0 32
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
44567.5 9
0
14 Logic Display~
6 1046 544 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44567.5 10
0
14 Logic Display~
6 995 546 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
44567.5 11
0
14 Logic Display~
6 954 552 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44567.5 12
0
14 Logic Display~
6 916 553 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44567.5 13
0
14 Logic Display~
6 869 556 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44567.5 14
0
14 Logic Display~
6 820 554 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
44567.5 15
0
14 Logic Display~
6 782 553 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
44567.5 16
0
14 Logic Display~
6 752 557 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
44567.5 17
0
14 Logic Display~
6 718 557 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
44567.5 18
0
14 Logic Display~
6 685 559 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
44567.5 19
0
14 Logic Display~
6 658 561 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
44567.5 20
0
4 4017
219 554 645 0 14 29
0 21 20 19 8 9 10 11 12 13
14 15 16 17 18
0
0 0 4832 0
4 4017
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 0 1 0 0 0
1 U
7678 0 0
2
44567.5 21
0
14 Logic Display~
6 789 274 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
44567.5 22
0
14 Logic Display~
6 758 269 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
44567.5 23
0
14 Logic Display~
6 731 262 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
44567.5 24
0
14 Logic Display~
6 701 261 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
44567.5 25
0
7 74LS569
162 528 284 0 18 37
0 7 6 5 32 31 30 29 28 27
26 4 3 33 2 25 24 23 22
0
0 0 4832 0
7 74LS569
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
162 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 9 7 12 2 1 11 6 5 4
3 8 17 18 19 13 14 15 16 9
7 12 2 1 11 6 5 4 3 8
17 18 19 13 14 15 16 0
65 0 0 512 1 0 0 0
1 U
8885 0 0
2
44567.5 26
0
31
1 14 2 0 0 8320 0 4 33 0 0 4
657 133
662 133
662 293
566 293
1 12 3 0 0 8320 0 5 33 0 0 4
601 149
606 149
606 258
566 258
1 11 4 0 0 8320 0 6 33 0 0 4
557 179
574 179
574 248
566 248
1 3 5 0 0 4224 0 1 33 0 0 4
315 233
472 233
472 266
490 266
1 2 6 0 0 4224 0 2 33 0 0 4
349 198
477 198
477 257
490 257
1 1 7 0 0 4224 0 3 33 0 0 4
296 171
482 171
482 248
490 248
4 1 8 0 0 4224 0 28 17 0 0 3
586 699
1046 699
1046 562
5 1 9 0 0 4224 0 28 18 0 0 3
586 690
995 690
995 564
6 1 10 0 0 4224 0 28 19 0 0 3
586 681
954 681
954 570
7 1 11 0 0 4224 0 28 20 0 0 3
586 672
916 672
916 571
8 1 12 0 0 4224 0 28 21 0 0 3
586 663
869 663
869 574
9 1 13 0 0 4224 0 28 22 0 0 3
586 654
820 654
820 572
10 1 14 0 0 4224 0 28 23 0 0 3
586 645
782 645
782 571
11 1 15 0 0 4224 0 28 24 0 0 3
586 636
752 636
752 575
12 1 16 0 0 4224 0 28 25 0 0 3
586 627
718 627
718 575
13 1 17 0 0 4224 0 28 26 0 0 3
586 618
685 618
685 577
14 1 18 0 0 4224 0 28 27 0 0 3
592 609
658 609
658 579
1 3 19 0 0 4224 0 7 28 0 0 4
411 707
508 707
508 690
522 690
1 2 20 0 0 4224 0 8 28 0 0 4
411 682
508 682
508 672
522 672
1 1 21 0 0 4224 0 9 28 0 0 4
412 657
508 657
508 663
516 663
18 1 22 0 0 4224 0 33 29 0 0 3
560 329
789 329
789 292
17 1 23 0 0 4224 0 33 30 0 0 3
560 320
758 320
758 287
16 1 24 0 0 4224 0 33 31 0 0 3
560 311
731 311
731 280
15 1 25 0 0 4224 0 33 32 0 0 3
560 302
701 302
701 279
1 10 26 0 0 4224 0 10 33 0 0 4
365 443
482 443
482 329
496 329
1 9 27 0 0 4224 0 11 33 0 0 4
366 416
467 416
467 320
496 320
1 8 28 0 0 4224 0 12 33 0 0 4
384 392
477 392
477 311
496 311
1 7 29 0 0 4224 0 13 33 0 0 4
359 347
472 347
472 302
496 302
1 6 30 0 0 4224 0 14 33 0 0 4
365 320
482 320
482 293
490 293
1 5 31 0 0 4224 0 15 33 0 0 4
424 304
477 304
477 284
496 284
1 4 32 0 0 4224 0 16 33 0 0 4
426 285
482 285
482 275
496 275
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
531 716 730 740
538 721 722 737
23 5-Stage Johnson Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
541 346 780 370
548 351 772 367
28 4-Bit Binary Up/Down Counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
