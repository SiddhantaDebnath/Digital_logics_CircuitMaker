CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
19 E:\Software\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
34
5 7415~
219 415 370 0 1 22
0 0
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
5130 0 0
2
44566.7 0
0
5 7415~
219 425 276 0 1 22
0 0
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
391 0 0
2
44566.7 0
0
5 7415~
219 421 180 0 1 22
0 0
0
0 0 608 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
3124 0 0
2
44566.7 0
0
13 Logic Switch~
5 344 514 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 782
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 235 507 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 782
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 149 506 0 1 11
0 11
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 349 1045 0 1 11
0 14
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 232 1045 0 1 11
0 13
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90014e-315 5.26354e-315
0
13 Logic Switch~
5 108 1056 0 1 11
0 12
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.90014e-315 5.30499e-315
0
13 Logic Switch~
5 263 60 0 1 11
0 28
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.90014e-315 5.36716e-315
0
13 Logic Switch~
5 167 60 0 1 11
0 30
0
0 0 21344 782
2 0V
-6 -20 8 -12
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.90014e-315 5.37752e-315
0
13 Logic Switch~
5 67 59 0 1 11
0 31
0
0 0 21344 782
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.90014e-315 5.38788e-315
0
5 7412~
219 654 669 0 4 22
0 5 4 3 2
0
0 0 608 0
4 7412
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 6 0
1 U
3536 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 819 631 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90014e-315 0
0
5 7412~
219 526 742 0 4 22
0 8 7 6 3
0
0 0 608 0
4 7412
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 5 0
1 U
3835 0 0
2
5.90014e-315 0
0
5 7412~
219 523 680 0 4 22
0 8 10 9 4
0
0 0 608 0
4 7412
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 5 0
1 U
3670 0 0
2
5.90014e-315 0
0
5 7412~
219 521 612 0 4 22
0 11 7 9 5
0
0 0 608 0
4 7412
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
5616 0 0
2
5.90014e-315 0
0
10 2-In NAND~
219 360 564 0 3 22
0 9 9 6
0
0 0 608 782
4 7400
-7 -24 21 -16
3 U4C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9323 0 0
2
5.90014e-315 0
0
10 2-In NAND~
219 255 560 0 3 22
0 10 10 7
0
0 0 608 782
4 7400
-7 -24 21 -16
3 U4B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
317 0 0
2
5.90014e-315 0
0
10 2-In NAND~
219 124 616 0 3 22
0 11 11 8
0
0 0 608 782
4 7400
-7 -24 21 -16
3 U4A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3108 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 940 1288 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44566.7 0
0
14 Logic Display~
6 747 264 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
44566.7 1
0
9 2-In NOR~
219 844 1318 0 3 22
0 20 20 19
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
7876 0 0
2
5.90014e-315 5.39306e-315
0
9 3-In NOR~
219 526 1444 0 4 22
0 12 13 14 21
0
0 0 608 0
6 74LS27
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 9 0
1 U
6369 0 0
2
5.90014e-315 5.39824e-315
0
9 3-In NOR~
219 713 1318 0 4 22
0 23 22 21 20
0
0 0 608 0
6 74LS27
-21 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 8 0
1 U
9172 0 0
2
5.90014e-315 5.40342e-315
0
9 3-In NOR~
219 525 1321 0 4 22
0 12 16 15 22
0
0 0 608 0
6 74LS27
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 8 0
1 U
7100 0 0
2
5.90014e-315 5.4086e-315
0
9 3-In NOR~
219 526 1228 0 4 22
0 17 13 15 23
0
0 0 608 0
6 74LS27
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 8 0
1 U
3820 0 0
2
5.90014e-315 5.41378e-315
0
9 2-In NOR~
219 395 1120 0 3 22
0 14 14 15
0
0 0 608 270
6 74LS02
-21 -24 21 -16
3 U7C
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
7678 0 0
2
5.90014e-315 5.41896e-315
0
9 2-In NOR~
219 277 1121 0 3 22
0 13 13 16
0
0 0 608 270
6 74LS02
-21 -24 21 -16
3 U7B
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
961 0 0
2
5.90014e-315 5.42414e-315
0
9 2-In NOR~
219 158 1112 0 3 22
0 12 12 17
0
0 0 608 270
6 74LS02
-21 -24 21 -16
3 U7A
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3178 0 0
2
5.90014e-315 5.42933e-315
0
8 3-In OR~
219 653 288 0 4 22
0 26 24 25 18
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
3409 0 0
2
5.90014e-315 5.45782e-315
0
9 Inverter~
13 300 108 0 2 22
0 28 27
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3951 0 0
2
5.90014e-315 5.46041e-315
0
9 Inverter~
13 205 109 0 2 22
0 30 29
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8885 0 0
2
5.90014e-315 5.463e-315
0
9 Inverter~
13 107 106 0 2 22
0 31 32
0
0 0 608 782
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3780 0 0
2
5.90014e-315 5.46559e-315
0
60
4 3 0 0 0 0 0 1 31 0 0 4
436 370
632 370
632 297
640 297
4 2 0 0 0 0 0 2 31 0 0 4
446 276
627 276
627 288
641 288
4 1 0 0 0 0 0 3 31 0 0 4
442 180
632 180
632 279
640 279
4 0 0 0 0 0 0 3 0 0 0 2
442 180
448 180
4 1 2 0 0 4224 0 13 14 0 0 3
681 669
819 669
819 649
4 3 3 0 0 4224 0 15 13 0 0 4
553 742
617 742
617 678
630 678
4 2 4 0 0 4224 0 16 13 0 0 4
550 680
622 680
622 669
630 669
4 1 5 0 0 4224 0 17 13 0 0 4
548 612
622 612
622 660
630 660
3 3 6 0 0 4224 0 18 15 0 0 3
361 590
361 751
502 751
0 2 7 0 0 4096 0 0 15 16 0 4
256 612
482 612
482 742
502 742
0 1 8 0 0 4096 0 0 15 14 0 4
125 671
494 671
494 733
502 733
0 3 9 0 0 12416 0 0 16 15 0 5
344 531
344 535
486 535
486 689
499 689
0 2 10 0 0 12416 0 0 16 21 0 4
235 526
330 526
330 680
499 680
3 1 8 0 0 8320 0 20 16 0 0 3
125 642
125 671
499 671
0 3 9 0 0 0 0 0 17 19 0 4
344 531
489 531
489 621
497 621
3 2 7 0 0 8320 0 19 17 0 0 3
256 586
256 612
497 612
0 1 11 0 0 4224 0 0 17 23 0 4
149 518
335 518
335 603
497 603
0 1 9 0 0 0 0 0 18 19 0 3
360 531
360 539
352 539
1 2 9 0 0 0 0 4 18 0 0 4
344 526
344 531
370 531
370 539
0 1 10 0 0 0 0 0 19 21 0 3
250 527
250 535
247 535
1 2 10 0 0 0 0 5 19 0 0 4
235 519
235 527
265 527
265 535
0 1 11 0 0 0 0 0 20 23 0 3
161 527
161 591
116 591
1 2 11 0 0 0 0 6 20 0 0 6
149 518
149 527
161 527
161 527
134 527
134 591
1 0 12 0 0 4096 0 9 0 0 45 2
108 1068
108 1080
1 0 13 0 0 4096 0 8 0 0 43 2
232 1057
232 1077
1 0 14 0 0 4096 0 7 0 0 41 2
349 1057
349 1076
0 2 13 0 0 8192 0 0 24 43 0 3
233 1228
233 1444
514 1444
0 1 12 0 0 8320 0 0 24 45 0 3
109 1312
109 1435
513 1435
0 3 15 0 0 4096 0 0 26 31 0 4
401 1235
504 1235
504 1330
512 1330
3 2 16 0 0 8320 0 29 26 0 0 3
283 1154
283 1321
513 1321
3 3 15 0 0 8320 0 28 27 0 0 3
401 1153
401 1237
513 1237
3 1 17 0 0 8320 0 30 27 0 0 3
164 1145
164 1219
513 1219
4 1 18 0 0 4224 0 31 22 0 0 3
686 288
747 288
747 282
3 1 19 0 0 4224 0 23 21 0 0 3
883 1318
940 1318
940 1306
0 2 20 0 0 8192 0 0 23 36 0 3
798 1318
798 1327
831 1327
4 1 20 0 0 4224 0 25 23 0 0 4
752 1318
798 1318
798 1309
831 1309
4 3 21 0 0 8320 0 24 25 0 0 4
565 1444
627 1444
627 1327
700 1327
4 2 22 0 0 12416 0 26 25 0 0 4
564 1321
627 1321
627 1318
701 1318
4 1 23 0 0 8320 0 27 25 0 0 4
565 1228
626 1228
626 1309
700 1309
0 1 14 0 0 0 0 0 28 41 0 3
392 1087
410 1087
410 1101
3 2 14 0 0 8320 0 24 28 0 0 5
513 1453
349 1453
349 1074
392 1074
392 1101
0 1 13 0 0 0 0 0 29 43 0 3
274 1086
292 1086
292 1102
2 2 13 0 0 4224 0 27 29 0 0 5
514 1228
232 1228
232 1072
274 1072
274 1102
1 2 12 0 0 0 0 30 30 0 0 2
173 1093
155 1093
1 2 12 0 0 0 0 26 30 0 0 5
512 1312
108 1312
108 1071
155 1071
155 1093
2 3 27 0 0 4224 0 32 1 0 0 5
303 126
303 380
394 380
394 379
391 379
1 1 28 0 0 8192 0 32 10 0 0 3
303 90
303 72
263 72
0 3 28 0 0 4096 0 0 3 49 0 2
263 189
397 189
0 0 28 0 0 0 0 0 0 0 50 2
391 189
263 189
1 3 28 0 0 4224 0 10 2 0 0 4
263 72
263 284
401 284
401 285
2 2 29 0 0 4224 0 33 1 0 0 5
208 127
208 371
394 371
394 370
391 370
0 2 30 0 0 8320 0 0 2 56 0 4
167 180
167 275
401 275
401 276
0 0 31 0 0 4096 0 0 0 59 0 2
67 170
67 173
0 2 29 0 0 0 0 0 33 0 0 2
208 130
208 127
1 1 30 0 0 0 0 11 33 0 0 3
167 72
208 72
208 91
1 2 30 0 0 0 0 11 3 0 0 3
167 72
167 180
397 180
0 1 32 0 0 16512 0 0 1 58 0 7
110 265
110 363
112 363
112 362
394 362
394 361
391 361
2 1 32 0 0 0 0 34 2 0 0 4
110 124
110 266
401 266
401 267
1 1 31 0 0 8320 0 12 3 0 0 3
67 71
67 171
397 171
1 1 31 0 0 0 0 12 34 0 0 4
67 71
67 76
110 76
110 88
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
746 1403 839 1427
756 1411 828 1427
9 NOR Logic
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
945 579 1046 603
955 587 1035 603
10 NAND Logic
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
820 102 913 126
830 110 902 126
9 AOI Logic
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
