CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
19 E:\Software\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 611 469 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -15 8 -7
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 603 374 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -15 8 -7
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 703 174 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.90014e-315 5.26354e-315
0
13 Logic Switch~
5 703 116 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 92 395 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.90014e-315 5.26354e-315
0
13 Logic Switch~
5 93 454 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 89 176 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.90014e-315 0
0
13 Logic Switch~
5 88 117 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 935 402 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 989 131 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 384 401 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.90014e-315 0
0
14 Logic Display~
6 351 116 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90014e-315 0
0
9 2-In AND~
219 232 419 0 3 22
0 16 15 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9265 0 0
2
5.90014e-315 0
0
9 Inverter~
13 799 175 0 2 22
0 12 10
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9442 0 0
2
5.90014e-315 5.30499e-315
0
9 2-In AND~
219 917 148 0 3 22
0 11 10 2
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9424 0 0
2
5.90014e-315 5.26354e-315
0
9 Inverter~
13 794 117 0 2 22
0 13 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
9968 0 0
2
5.90014e-315 0
0
9 Inverter~
13 318 419 0 2 22
0 14 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
9281 0 0
2
5.90014e-315 0
0
9 Inverter~
13 702 469 0 2 22
0 8 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
8464 0 0
2
5.90014e-315 0
0
9 Inverter~
13 696 373 0 2 22
0 9 7
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
7168 0 0
2
5.90014e-315 0
0
9 Inverter~
13 284 147 0 2 22
0 17 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3171 0 0
2
5.90014e-315 0
0
8 2-In OR~
219 844 421 0 3 22
0 7 6 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4139 0 0
2
5.90014e-315 0
0
8 2-In OR~
219 204 147 0 3 22
0 19 18 17
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6435 0 0
2
5.90014e-315 0
0
18
3 1 2 0 0 4224 0 15 10 0 0 4
938 148
974 148
974 149
989 149
3 1 3 0 0 8320 0 21 9 0 0 3
877 421
877 420
935 420
2 1 4 0 0 4224 0 17 11 0 0 2
339 419
384 419
2 1 5 0 0 4224 0 20 12 0 0 3
305 147
351 147
351 134
2 2 6 0 0 4224 0 18 21 0 0 4
723 469
793 469
793 430
831 430
2 1 7 0 0 4224 0 19 21 0 0 4
717 373
792 373
792 412
831 412
1 1 8 0 0 4224 0 1 18 0 0 2
623 469
687 469
1 1 9 0 0 8320 0 2 19 0 0 3
615 374
615 373
681 373
2 2 10 0 0 8320 0 14 15 0 0 3
820 175
820 157
893 157
2 1 11 0 0 8320 0 16 15 0 0 3
815 117
815 139
893 139
1 1 12 0 0 4224 0 3 14 0 0 4
715 174
769 174
769 175
784 175
1 1 13 0 0 8320 0 4 16 0 0 3
715 116
715 117
779 117
3 1 14 0 0 4224 0 13 17 0 0 2
253 419
303 419
1 2 15 0 0 12416 0 6 13 0 0 4
105 454
152 454
152 428
208 428
1 1 16 0 0 12416 0 5 13 0 0 4
104 395
152 395
152 410
208 410
3 1 17 0 0 4224 0 22 20 0 0 2
237 147
269 147
1 2 18 0 0 8320 0 7 22 0 0 3
101 176
101 156
191 156
1 1 19 0 0 8320 0 8 22 0 0 3
100 117
100 138
191 138
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
77 61 138 85
87 69 127 85
5 LHS:-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
694 48 755 72
704 56 744 72
5 RHS:-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
594 321 655 345
604 329 644 345
5 RHS:-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
64 342 125 366
74 350 114 366
5 LHS:-
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
78 278 147 302
88 286 136 302
6 Law 2:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
56 0 125 24
66 8 114 24
6 Law 1:
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
